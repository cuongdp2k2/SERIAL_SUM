module Hex_to_Dec (
    // input 
        input logic [1:0][7:0] Hex_i ,

    // output
        output logic            Carry_o ,
        output logic [2:0][7:0] Dec_o 
);
endmodule : Hex_to_Dec
